//-----------------------------------------------------
// File Name   : alucodes.sv
// Function    : pMIPS ALU function code definitions 
//-----------------------------------------------------
// 
`define RADD  1'b0
`define RMUL  1'b1   // new multiply

